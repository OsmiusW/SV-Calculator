`timescale 1ns/1ps

module InstructionSet
	#(parameter WIDTH = 32)
	(input logic [WIDTH-1:0] Instruction,
	output logic [WIDTH-1:0] Set);
	
	
assign 	
	
endmodule