`timescale 1ns / 1ps

module Controller 
	input logic [6:0] OpCode,
	output logic [3:0] ALU,
	output logic MEM,
	output logic ImmValue,
	output logic RegValue,
	
	assign MEM = ;
	assign ImmValue = ;
	assign RegValue = ;
	
endmodule